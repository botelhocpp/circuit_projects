CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 60 10
133 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
301 176 414 273
42991634 0
0
6 Title:
5 Name:
0
0
0
62
13 Logic Switch~
5 45 414 0 1 11
0 23
0
0 0 21872 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
5 CLOCK
-16 -32 19 -24
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3795 0 0
2
45461.7 0
0
13 Logic Switch~
5 44 475 0 1 11
0 24
0
0 0 21872 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
5 RESET
-17 -31 18 -23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3637 0 0
2
45461.7 1
0
13 Logic Switch~
5 48 314 0 1 11
0 100
0
0 0 21872 0
2 0V
-7 -17 7 -9
2 V2
-6 -26 8 -18
4 Inic
-13 -30 15 -22
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3226 0 0
2
45461.7 2
0
12 Hex Display~
7 1461 353 0 16 19
10 14 13 12 11 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP7
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6966 0 0
2
45461.7 3
0
12 Hex Display~
7 1497 353 0 16 19
10 18 17 16 15 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP6
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9796 0 0
2
45461.7 4
0
14 Logic Display~
6 2080 812 0 1 2
10 21
0
0 0 54384 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
3 FIM
-11 -23 10 -15
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5952 0 0
2
45461.7 5
0
7 Ground~
168 1948 815 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3649 0 0
2
45461.7 6
0
5 4071~
219 1876 845 0 3 22
0 27 26 22
0
0 0 1136 0
4 4071
-7 -24 21 -16
3 U4D
-3 -25 18 -17
5 �LOAD
-10 -28 25 -20
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
3716 0 0
2
45461.7 7
0
5 4049~
219 1821 875 0 2 22
0 25 26
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 5 0
1 U
4797 0 0
2
45461.7 8
0
5 4081~
219 1711 836 0 3 22
0 29 28 27
0
0 0 1136 0
4 4081
-7 -24 21 -16
4 U22A
-15 -25 13 -17
4 �R/W
-17 -29 11 -21
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
4681 0 0
2
45461.7 9
0
5 4013~
219 1970 881 0 6 22
0 2 22 23 24 105 21
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U21A
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 7 0
1 U
9730 0 0
2
45461.7 10
0
7 Ground~
168 1583 998 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9874 0 0
2
45461.7 11
0
2 +V
167 1594 695 0 1 3
0 30
0
0 0 54256 0
2 5V
-9 -22 5 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
364 0 0
2
45461.7 12
0
4 4585
219 1638 906 0 14 29
0 15 16 17 18 30 30 30 30 2
30 2 106 28 107
0
0 0 4848 0
4 4585
-14 -60 14 -52
3 U20
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
3656 0 0
2
45461.7 13
0
4 4585
219 1637 757 0 14 29
0 11 12 13 14 30 30 30 30 2
30 2 108 29 109
0
0 0 4848 0
4 4585
-14 -60 14 -52
3 U19
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
3131 0 0
2
45461.7 14
0
7 Ground~
168 1340 587 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6772 0 0
2
45461.7 15
0
4 4076
219 1815 591 0 22 29
0 43 42 41 40 19 19 31 31 23
24 39 38 37 36 0 0 0 0 0
0 0 1
0
0 0 4848 0
4 4076
-14 -60 14 -52
3 U18
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 14 10 9 2 1 7
15 3 4 5 6 11 12 13 14 10
9 2 1 7 15 3 4 5 6 0
65 0 0 0 1 0 0 0
1 U
9557 0 0
2
45461.7 16
0
4 4076
219 1816 444 0 14 29
0 47 46 45 44 19 19 31 31 23
24 35 34 33 32
0
0 0 4848 0
4 4076
-14 -60 14 -52
3 U17
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 14 10 9 2 1 7
15 3 4 5 6 11 12 13 14 10
9 2 1 7 15 3 4 5 6 0
65 0 0 0 1 0 0 0
1 U
5789 0 0
2
45461.7 17
0
7 74LS244
143 1642 597 0 18 37
0 32 33 34 35 36 37 38 39 11
12 13 14 15 16 17 18 31 31
0
0 0 4848 512
7 74LS244
-24 -60 25 -52
3 U16
-17 -61 4 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 0 0 0
1 U
7328 0 0
2
45461.7 18
0
7 74LS244
143 1637 435 0 18 37
0 11 12 13 14 15 16 17 18 47
46 45 44 43 42 41 40 19 19
0
0 0 4848 0
7 74LS244
-24 -60 25 -52
3 U15
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP14
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 0 0 0
1 U
4799 0 0
2
45461.7 19
0
5 4049~
219 1425 248 0 2 22
0 19 31
0
0 0 624 270
4 4049
-7 -24 21 -16
3 U5C
16 -8 37 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 5 0
1 U
9196 0 0
2
45461.7 20
0
6 1K RAM
79 1382 426 0 20 41
0 2 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 64
31
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
3 U14
-11 -70 10 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 0 1 0 0 0
1 U
3857 0 0
2
45461.7 21
0
7 Ground~
168 1189 584 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7125 0 0
2
45461.7 22
0
7 74LS157
122 1233 517 0 14 29
0 19 52 59 53 58 54 57 55 56
2 3 4 5 6
0
0 0 4848 0
7 74F157A
-24 -60 25 -52
3 U12
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3641 0 0
2
45461.7 23
0
7 74LS157
122 1237 348 0 14 29
0 19 48 63 49 62 50 61 51 60
2 7 8 9 10
0
0 0 4848 0
7 74F157A
-24 -60 25 -52
3 U13
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
9821 0 0
2
45461.7 24
0
2 +V
167 828 184 0 1 3
0 65
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3187 0 0
2
45461.7 25
0
14 Logic Display~
6 657 154 0 1 2
10 64
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
762 0 0
2
45461.7 26
0
14 Logic Display~
6 637 154 0 1 2
10 66
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
39 0 0
2
45461.7 27
0
14 Logic Display~
6 614 155 0 1 2
10 67
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9450 0 0
2
45461.7 28
0
14 Logic Display~
6 592 155 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3236 0 0
2
5.90128e-315 0
0
14 Logic Display~
6 448 153 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3321 0 0
2
5.90128e-315 5.26354e-315
0
14 Logic Display~
6 426 153 0 1 2
10 68
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8879 0 0
2
5.90128e-315 5.30499e-315
0
12 Hex Display~
7 983 839 0 16 19
10 69 70 71 72 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP5
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5433 0 0
2
5.90128e-315 5.32571e-315
0
12 Hex Display~
7 970 490 0 18 19
10 55 54 53 52 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3679 0 0
2
5.90128e-315 5.34643e-315
0
12 Hex Display~
7 1010 490 0 18 19
10 51 50 49 48 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9342 0 0
2
5.90128e-315 5.3568e-315
0
12 Hex Display~
7 971 245 0 18 19
10 56 57 58 59 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3623 0 0
2
5.90128e-315 5.36716e-315
0
12 Hex Display~
7 1008 245 0 18 19
10 60 61 62 63 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3722 0 0
2
5.90128e-315 5.37752e-315
0
8 Hex Key~
166 149 832 0 11 12
0 74 75 76 77 0 0 0 0 0
4 52
0
0 0 4656 0
0
4 KPD5
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8993 0 0
2
5.90128e-315 5.38788e-315
0
8 Hex Key~
166 112 687 0 11 12
0 78 79 80 81 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD4
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3723 0 0
2
5.90128e-315 5.39306e-315
0
8 Hex Key~
166 149 687 0 11 12
0 82 83 84 85 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6244 0 0
2
5.90128e-315 5.39824e-315
0
7 74LS193
137 902 860 0 14 29
0 65 66 67 24 77 76 75 74 110
25 72 71 70 69
0
0 0 4848 0
6 74F193
-21 -51 21 -43
3 U11
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
6421 0 0
2
5.90128e-315 5.40342e-315
0
7 74LS193
137 894 637 0 14 29
0 73 65 67 24 81 80 79 78 111
112 52 53 54 55
0
0 0 4848 0
6 74F193
-21 -51 21 -43
3 U10
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
7743 0 0
2
5.90128e-315 5.4086e-315
0
7 74LS193
137 894 514 0 14 29
0 66 65 67 24 85 84 83 82 73
113 48 49 50 51
0
0 0 4848 0
6 74F193
-21 -51 21 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9840 0 0
2
5.90128e-315 5.41378e-315
0
8 Hex Key~
166 147 551 0 11 12
0 90 91 92 93 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6910 0 0
2
5.90128e-315 5.41896e-315
0
8 Hex Key~
166 110 550 0 11 12
0 86 87 88 89 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
449 0 0
2
5.90128e-315 5.42414e-315
0
7 74LS193
137 895 390 0 14 29
0 94 65 67 24 89 88 87 86 114
115 59 58 57 56
0
0 0 4848 0
6 74F193
-21 -51 21 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
8761 0 0
2
5.90128e-315 5.42933e-315
0
7 74LS193
137 895 269 0 14 29
0 66 65 67 24 93 92 91 90 94
116 63 62 61 60
0
0 0 4848 0
6 74F193
-21 -51 21 -43
2 U7
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
6748 0 0
2
5.90128e-315 5.43192e-315
0
5 4081~
219 190 224 0 3 22
0 68 95 97
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
7393 0 0
2
5.90128e-315 5.43451e-315
0
5 4071~
219 245 195 0 3 22
0 98 97 96
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
7699 0 0
2
5.90128e-315 5.4371e-315
0
7 Ground~
168 306 312 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6638 0 0
2
5.90128e-315 5.43969e-315
0
7 Ground~
168 306 164 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4595 0 0
2
5.90128e-315 5.44228e-315
0
10 2-In XNOR~
219 541 371 0 3 22
0 68 20 64
0
0 0 1136 0
4 4077
-7 -24 21 -16
3 U6A
-5 -25 16 -17
3 �CE
-7 -26 14 -18
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
9395 0 0
2
45461.7 29
0
5 4071~
219 540 260 0 3 22
0 68 20 67
0
0 0 1136 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
5 �LOAD
-10 -28 25 -20
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
3303 0 0
2
45461.7 30
0
5 4081~
219 548 315 0 3 22
0 68 20 66
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U3C
-12 -25 9 -17
5 COUNT
-18 -27 17 -19
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
4498 0 0
2
45461.7 31
0
5 4081~
219 548 204 0 3 22
0 68 95 19
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
4 �R/W
-17 -29 11 -21
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
9728 0 0
2
45461.7 32
0
5 4049~
219 102 177 0 2 22
0 22 103
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
3789 0 0
2
45461.7 33
0
5 4049~
219 97 314 0 2 22
0 100 99
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
3978 0 0
2
45461.7 34
0
5 4071~
219 243 341 0 3 22
0 104 68 101
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3494 0 0
2
45461.7 35
0
5 4081~
219 196 305 0 3 22
0 95 99 104
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3507 0 0
2
45461.7 36
0
9 3-In AND~
219 188 168 0 4 22
0 20 102 103 98
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 2 0
1 U
5151 0 0
2
45461.7 37
0
5 4013~
219 322 377 0 6 22
0 2 101 23 24 95 20
0
0 0 5744 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
2 Q0
5 7 19 15
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 2 1 0
1 U
3701 0 0
2
45461.7 38
0
5 4013~
219 321 231 0 6 22
0 2 96 23 24 102 68
0
0 0 5744 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
2 Q1
7 3 21 11
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 1 0
1 U
8585 0 0
2
45461.7 39
0
216
11 3 3 0 0 8320 0 24 22 0 0 4
1265 499
1294 499
1294 408
1350 408
4 12 4 0 0 8320 0 22 24 0 0 4
1350 417
1299 417
1299 517
1265 517
13 5 5 0 0 8320 0 24 22 0 0 4
1265 535
1305 535
1305 426
1350 426
14 6 6 0 0 8320 0 24 22 0 0 4
1265 553
1310 553
1310 435
1350 435
7 11 7 0 0 8320 0 22 25 0 0 4
1350 444
1315 444
1315 330
1269 330
8 12 8 0 0 8320 0 22 25 0 0 4
1350 453
1322 453
1322 348
1269 348
13 9 9 0 0 8320 0 25 22 0 0 4
1269 366
1327 366
1327 462
1350 462
14 10 10 0 0 8320 0 25 22 0 0 4
1269 384
1333 384
1333 471
1350 471
4 0 11 0 0 4096 0 4 0 0 100 2
1452 377
1452 408
3 0 12 0 0 4096 0 4 0 0 99 2
1458 377
1458 417
2 0 13 0 0 4096 0 4 0 0 98 2
1464 377
1464 426
1 0 14 0 0 4096 0 4 0 0 97 2
1470 377
1470 435
4 0 15 0 0 4096 0 5 0 0 95 2
1488 377
1488 444
3 0 16 0 0 4096 0 5 0 0 94 2
1494 377
1494 453
2 0 17 0 0 4096 0 5 0 0 93 2
1500 377
1500 462
1 0 18 0 0 4096 0 5 0 0 92 2
1506 377
1506 471
1 0 19 0 0 4096 0 21 0 0 82 2
1428 230
1428 205
1 0 20 0 0 4096 0 31 0 0 205 2
448 171
448 269
6 1 21 0 0 4224 0 11 6 0 0 3
1994 845
2080 845
2080 830
1 1 2 0 0 4096 0 11 7 0 0 4
1970 824
1970 789
1948 789
1948 809
1 0 22 0 0 12416 0 56 0 0 28 5
87 177
60 177
60 66
1921 66
1921 845
0 0 23 0 0 4096 0 0 0 75 25 2
1766 636
1766 1033
0 0 24 0 0 4096 0 0 0 80 24 2
1771 645
1771 1047
4 0 24 0 0 8320 0 11 0 0 211 4
1970 887
1970 1047
73 1047
73 475
0 3 23 0 0 8320 0 0 11 208 0 5
84 414
84 1033
1919 1033
1919 863
1946 863
1 10 25 0 0 12416 0 9 41 0 0 6
1806 875
1691 875
1691 1020
955 1020
955 860
940 860
2 2 26 0 0 8320 0 8 9 0 0 4
1863 854
1853 854
1853 875
1842 875
3 2 22 0 0 0 0 8 11 0 0 2
1909 845
1946 845
3 1 27 0 0 4224 0 10 8 0 0 2
1732 836
1863 836
2 13 28 0 0 8320 0 10 14 0 0 4
1687 845
1682 845
1682 915
1670 915
13 1 29 0 0 8320 0 15 10 0 0 4
1669 766
1680 766
1680 827
1687 827
1 0 30 0 0 4096 0 13 0 0 45 2
1594 704
1594 757
0 1 2 0 0 0 0 0 12 35 0 3
1584 969
1583 969
1583 992
9 0 2 0 0 0 0 14 0 0 35 2
1606 951
1584 951
11 0 2 0 0 8192 0 14 0 0 36 3
1606 969
1584 969
1584 820
9 11 2 0 0 0 0 15 15 0 0 4
1605 802
1584 802
1584 820
1605 820
6 0 30 0 0 0 0 14 0 0 40 2
1606 915
1593 915
7 0 30 0 0 0 0 14 0 0 40 2
1606 924
1593 924
10 0 30 0 0 0 0 14 0 0 40 3
1606 960
1594 960
1594 933
8 0 30 0 0 0 0 14 0 0 41 3
1606 933
1593 933
1593 906
0 5 30 0 0 4224 0 0 14 42 0 3
1593 811
1593 906
1606 906
10 0 30 0 0 0 0 15 0 0 45 3
1605 811
1593 811
1593 784
0 6 30 0 0 0 0 0 15 45 0 3
1593 767
1593 766
1605 766
7 0 30 0 0 0 0 15 0 0 45 2
1605 775
1593 775
5 8 30 0 0 0 0 15 15 0 0 4
1605 757
1593 757
1593 784
1605 784
4 0 18 0 0 8320 0 14 0 0 85 3
1606 897
1527 897
1527 642
3 0 17 0 0 8320 0 14 0 0 86 3
1606 888
1533 888
1533 633
2 0 16 0 0 8320 0 14 0 0 87 3
1606 879
1538 879
1538 624
1 0 15 0 0 8320 0 14 0 0 88 3
1606 870
1543 870
1543 615
4 0 14 0 0 8192 0 15 0 0 89 3
1605 748
1548 748
1548 597
0 3 13 0 0 4096 0 0 15 90 0 3
1555 588
1555 739
1605 739
2 0 12 0 0 8192 0 15 0 0 91 3
1605 730
1561 730
1561 579
1 0 11 0 0 8192 0 15 0 0 84 3
1605 721
1568 721
1568 570
0 1 2 0 0 4096 0 0 16 119 0 2
1340 398
1340 581
0 0 31 0 0 8192 0 0 0 79 81 4
1761 627
1725 627
1725 532
1682 532
0 0 19 0 0 12288 0 0 0 76 96 5
1756 609
1730 609
1730 495
1595 495
1595 444
1 14 32 0 0 16512 0 19 18 0 0 6
1668 570
1707 570
1707 695
1897 695
1897 408
1848 408
13 2 33 0 0 8320 0 18 19 0 0 6
1848 417
1891 417
1891 690
1702 690
1702 579
1668 579
3 12 34 0 0 16512 0 19 18 0 0 6
1668 588
1698 588
1698 685
1885 685
1885 426
1848 426
4 11 35 0 0 16512 0 19 18 0 0 6
1668 597
1693 597
1693 680
1879 680
1879 435
1848 435
14 5 36 0 0 12416 0 17 19 0 0 6
1847 555
1874 555
1874 675
1688 675
1688 615
1668 615
13 6 37 0 0 12416 0 17 19 0 0 6
1847 564
1868 564
1868 671
1684 671
1684 624
1668 624
12 7 38 0 0 12416 0 17 19 0 0 6
1847 573
1862 573
1862 666
1679 666
1679 633
1668 633
11 8 39 0 0 12416 0 17 19 0 0 6
1847 582
1856 582
1856 661
1674 661
1674 642
1668 642
4 16 40 0 0 8320 0 17 20 0 0 4
1783 582
1736 582
1736 480
1669 480
15 3 41 0 0 8320 0 20 17 0 0 4
1669 471
1740 471
1740 573
1783 573
2 14 42 0 0 8320 0 17 20 0 0 4
1783 564
1745 564
1745 462
1669 462
13 1 43 0 0 8320 0 20 17 0 0 4
1669 453
1751 453
1751 555
1783 555
4 12 44 0 0 4224 0 18 20 0 0 2
1784 435
1669 435
11 3 45 0 0 4224 0 20 18 0 0 2
1669 426
1784 426
2 10 46 0 0 4224 0 18 20 0 0 2
1784 417
1669 417
0 0 19 0 0 4096 0 0 0 76 77 2
1756 600
1756 460
0 0 31 0 0 4096 0 0 0 78 79 2
1761 479
1761 618
9 1 47 0 0 4224 0 20 18 0 0 2
1669 408
1784 408
9 9 23 0 0 0 0 18 17 0 0 4
1784 489
1766 489
1766 636
1783 636
5 6 19 0 0 0 0 17 17 0 0 4
1777 600
1756 600
1756 609
1777 609
5 6 19 0 0 0 0 18 18 0 0 4
1778 453
1756 453
1756 462
1778 462
7 8 31 0 0 0 0 18 18 0 0 4
1778 471
1761 471
1761 480
1778 480
7 8 31 0 0 0 0 17 17 0 0 4
1777 618
1761 618
1761 627
1777 627
10 10 24 0 0 0 0 18 17 0 0 4
1784 498
1771 498
1771 645
1783 645
0 0 31 0 0 4224 0 0 0 118 83 5
1428 399
1575 399
1575 532
1682 532
1682 561
0 0 19 0 0 8192 0 0 0 120 96 4
1181 204
1181 205
1595 205
1595 399
17 18 31 0 0 0 0 19 19 0 0 4
1674 561
1682 561
1682 606
1674 606
9 0 11 0 0 8192 0 19 0 0 100 3
1604 570
1567 570
1567 408
16 0 18 0 0 0 0 19 0 0 92 3
1604 642
1526 642
1526 471
15 0 17 0 0 0 0 19 0 0 93 3
1604 633
1533 633
1533 462
14 0 16 0 0 0 0 19 0 0 94 3
1604 624
1538 624
1538 453
13 0 15 0 0 0 0 19 0 0 95 3
1604 615
1543 615
1543 444
12 0 14 0 0 8192 0 19 0 0 97 3
1604 597
1548 597
1548 435
11 0 13 0 0 8192 0 19 0 0 98 3
1604 588
1554 588
1554 426
10 0 12 0 0 8192 0 19 0 0 99 3
1604 579
1561 579
1561 417
18 8 18 0 0 0 0 22 20 0 0 4
1414 471
1581 471
1581 480
1605 480
7 17 17 0 0 0 0 20 22 0 0 4
1605 471
1584 471
1584 462
1414 462
16 6 16 0 0 0 0 22 20 0 0 4
1414 453
1588 453
1588 462
1605 462
5 15 15 0 0 0 0 20 22 0 0 4
1605 453
1591 453
1591 444
1414 444
17 18 19 0 0 0 0 20 20 0 0 4
1599 399
1595 399
1595 444
1599 444
14 4 14 0 0 4224 0 22 20 0 0 2
1414 435
1605 435
3 13 13 0 0 4224 0 20 22 0 0 2
1605 426
1414 426
12 2 12 0 0 4224 0 22 20 0 0 2
1414 417
1605 417
11 1 11 0 0 4224 0 22 20 0 0 2
1414 408
1605 408
0 2 48 0 0 8320 0 0 25 139 0 4
1001 523
1108 523
1108 321
1205 321
0 4 49 0 0 8320 0 0 25 140 0 4
1007 532
1115 532
1115 339
1205 339
6 0 50 0 0 8320 0 25 0 0 141 4
1205 357
1120 357
1120 541
1013 541
0 8 51 0 0 8320 0 0 25 142 0 4
1018 550
1125 550
1125 375
1205 375
2 0 52 0 0 12416 0 24 0 0 146 4
1201 490
1131 490
1131 646
961 646
0 4 53 0 0 4224 0 0 24 145 0 4
966 655
1137 655
1137 508
1201 508
6 0 54 0 0 12416 0 24 0 0 144 4
1201 526
1143 526
1143 664
973 664
0 8 55 0 0 4224 0 0 24 143 0 4
979 673
1149 673
1149 544
1201 544
9 0 56 0 0 12416 0 24 0 0 135 4
1201 553
1157 553
1157 426
979 426
7 0 57 0 0 12416 0 24 0 0 136 4
1201 535
1162 535
1162 417
974 417
5 0 58 0 0 12416 0 24 0 0 137 4
1201 517
1169 517
1169 408
967 408
3 0 59 0 0 12416 0 24 0 0 138 4
1201 499
1175 499
1175 398
962 398
9 0 60 0 0 12416 0 25 0 0 132 4
1205 384
1159 384
1159 305
1017 305
0 7 61 0 0 4224 0 0 25 124 0 4
1011 295
1165 295
1165 366
1205 366
5 0 62 0 0 12416 0 25 0 0 133 4
1205 348
1171 348
1171 287
1004 287
0 3 63 0 0 4224 0 0 25 134 0 4
999 277
1176 277
1176 330
1205 330
0 19 64 0 0 8320 0 0 22 126 0 5
657 369
657 795
1436 795
1436 390
1420 390
2 20 31 0 0 0 0 21 22 0 0 3
1428 266
1428 399
1420 399
1 2 2 0 0 0 0 22 22 0 0 4
1350 390
1340 390
1340 399
1350 399
0 0 19 0 0 4224 0 0 0 129 123 3
592 204
1182 204
1182 312
10 0 2 0 0 0 0 24 0 0 122 2
1195 562
1189 562
10 1 2 0 0 8320 0 25 23 0 0 3
1199 393
1189 393
1189 578
1 1 19 0 0 0 0 25 24 0 0 4
1205 312
1182 312
1182 481
1201 481
2 13 61 0 0 0 0 37 47 0 0 5
1011 269
1011 295
1012 295
1012 296
927 296
0 1 65 0 0 4096 0 0 26 156 0 2
828 252
828 193
1 3 64 0 0 0 0 27 52 0 0 3
657 172
657 371
580 371
1 0 66 0 0 4096 0 28 0 0 187 2
637 172
637 315
1 0 67 0 0 4096 0 29 0 0 131 2
614 173
614 260
3 1 19 0 0 0 0 55 30 0 0 3
569 204
592 204
592 173
1 0 68 0 0 4096 0 32 0 0 207 2
426 171
426 195
0 3 67 0 0 4224 0 0 53 162 0 2
837 260
573 260
14 1 60 0 0 0 0 47 37 0 0 3
927 305
1017 305
1017 269
12 3 62 0 0 0 0 47 37 0 0 3
927 287
1005 287
1005 269
4 11 63 0 0 0 0 37 47 0 0 5
999 269
999 277
1000 277
1000 278
927 278
14 1 56 0 0 0 0 46 36 0 0 3
927 426
980 426
980 269
2 13 57 0 0 0 0 36 46 0 0 3
974 269
974 417
927 417
12 3 58 0 0 0 0 46 36 0 0 3
927 408
968 408
968 269
4 11 59 0 0 0 0 36 46 0 0 5
962 269
962 398
961 398
961 399
927 399
4 11 48 0 0 0 0 35 43 0 0 3
1001 514
1001 523
926 523
12 3 49 0 0 0 0 43 35 0 0 3
926 532
1007 532
1007 514
2 13 50 0 0 0 0 35 43 0 0 3
1013 514
1013 541
926 541
14 1 51 0 0 0 0 43 35 0 0 3
926 550
1019 550
1019 514
14 1 55 0 0 0 0 42 34 0 0 3
926 673
979 673
979 514
2 13 54 0 0 0 0 34 42 0 0 3
973 514
973 664
926 664
12 3 53 0 0 0 0 42 34 0 0 3
926 655
967 655
967 514
4 11 52 0 0 0 0 34 42 0 0 3
961 514
961 646
926 646
1 14 69 0 0 8320 0 33 41 0 0 3
992 863
992 896
934 896
13 2 70 0 0 4224 0 41 33 0 0 3
934 887
986 887
986 863
3 12 71 0 0 8320 0 33 41 0 0 3
980 863
980 878
934 878
11 4 72 0 0 4224 0 41 33 0 0 3
934 869
974 869
974 863
2 0 66 0 0 8320 0 41 0 0 155 3
870 842
821 842
821 487
0 1 65 0 0 4224 0 0 41 158 0 3
830 619
830 833
870 833
3 0 67 0 0 0 0 41 0 0 159 3
864 851
837 851
837 628
0 4 24 0 0 0 0 0 41 164 0 3
843 637
843 860
870 860
1 0 66 0 0 0 0 43 0 0 187 3
862 487
821 487
821 242
0 2 65 0 0 0 0 0 47 157 0 3
828 373
828 251
863 251
0 2 65 0 0 0 0 0 46 158 0 3
828 497
828 372
863 372
2 2 65 0 0 0 0 42 43 0 0 4
862 619
828 619
828 496
862 496
0 3 67 0 0 0 0 0 42 161 0 3
837 504
837 628
856 628
4 0 24 0 0 0 0 43 0 0 164 2
862 514
843 514
0 3 67 0 0 0 0 0 43 162 0 3
837 380
837 505
856 505
3 3 67 0 0 0 0 47 46 0 0 4
857 260
837 260
837 381
857 381
0 4 24 0 0 0 0 0 47 164 0 3
843 392
843 269
863 269
4 4 24 0 0 0 0 42 46 0 0 4
862 637
843 637
843 390
863 390
9 1 73 0 0 12416 0 43 42 0 0 6
932 505
943 505
943 574
849 574
849 610
862 610
8 1 74 0 0 4224 0 41 38 0 0 3
870 896
158 896
158 856
7 2 75 0 0 4224 0 41 38 0 0 3
870 887
152 887
152 856
3 6 76 0 0 8320 0 38 41 0 0 3
146 856
146 878
870 878
5 4 77 0 0 4224 0 41 38 0 0 3
870 869
140 869
140 856
8 1 78 0 0 12416 0 42 39 0 0 5
862 673
808 673
808 785
121 785
121 711
2 7 79 0 0 8320 0 39 42 0 0 5
115 711
115 775
799 775
799 664
862 664
6 3 80 0 0 12416 0 42 39 0 0 5
862 655
791 655
791 764
109 764
109 711
4 5 81 0 0 8320 0 39 42 0 0 5
103 711
103 753
784 753
784 646
862 646
8 1 82 0 0 12416 0 43 40 0 0 5
862 550
777 550
777 747
158 747
158 711
2 7 83 0 0 8320 0 40 43 0 0 5
152 711
152 739
769 739
769 541
862 541
6 3 84 0 0 12416 0 43 40 0 0 5
862 532
762 532
762 730
146 730
146 711
4 5 85 0 0 8320 0 40 43 0 0 5
140 711
140 721
753 721
753 523
862 523
8 1 86 0 0 12416 0 46 45 0 0 5
863 426
745 426
745 642
119 642
119 574
2 7 87 0 0 8320 0 45 46 0 0 5
113 574
113 632
733 632
733 417
863 417
6 3 88 0 0 12416 0 46 45 0 0 5
863 408
723 408
723 624
107 624
107 574
5 4 89 0 0 12416 0 46 45 0 0 5
863 399
714 399
714 616
101 616
101 574
1 8 90 0 0 8320 0 44 47 0 0 5
156 575
156 607
706 607
706 305
863 305
7 2 91 0 0 12416 0 47 44 0 0 5
863 296
698 296
698 598
150 598
150 575
3 6 92 0 0 8320 0 44 47 0 0 5
144 575
144 591
690 591
690 287
863 287
5 4 93 0 0 12416 0 47 44 0 0 5
863 278
683 278
683 583
138 583
138 575
0 0 24 0 0 0 0 0 0 211 163 4
281 475
675 475
675 269
843 269
3 1 66 0 0 0 0 54 47 0 0 4
569 315
668 315
668 242
863 242
9 1 94 0 0 12416 0 47 46 0 0 6
933 260
943 260
943 328
848 328
848 363
863 363
2 0 95 0 0 4096 0 48 0 0 197 2
166 233
148 233
0 1 20 0 0 8320 0 0 60 205 0 5
384 269
384 87
157 87
157 159
164 159
3 2 96 0 0 4224 0 49 62 0 0 2
278 195
297 195
1 0 68 0 0 4096 0 48 0 0 196 2
166 215
126 215
2 3 97 0 0 8320 0 49 48 0 0 4
232 204
220 204
220 224
211 224
4 1 98 0 0 8320 0 60 49 0 0 4
209 168
220 168
220 186
232 186
2 2 99 0 0 4224 0 59 57 0 0 2
172 314
118 314
0 2 68 0 0 12416 0 0 58 207 0 5
364 195
364 107
126 107
126 350
230 350
0 1 95 0 0 8320 0 0 59 206 0 5
394 215
394 79
148 79
148 296
172 296
1 1 2 0 0 0 0 50 61 0 0 4
306 306
306 296
322 296
322 320
1 1 2 0 0 0 0 62 51 0 0 4
321 174
321 148
306 148
306 158
2 0 20 0 0 0 0 54 0 0 202 2
524 324
487 324
1 0 68 0 0 0 0 53 0 0 204 2
527 251
503 251
0 2 20 0 0 0 0 0 52 205 0 3
487 269
487 380
525 380
0 1 68 0 0 0 0 0 52 204 0 3
503 306
503 362
525 362
0 1 68 0 0 0 0 0 54 207 0 3
503 195
503 306
524 306
2 6 20 0 0 0 0 53 61 0 0 4
527 269
384 269
384 341
346 341
5 2 95 0 0 0 0 61 55 0 0 4
352 359
394 359
394 213
524 213
6 1 68 0 0 0 0 62 55 0 0 2
345 195
524 195
0 1 23 0 0 0 0 0 1 209 0 3
291 359
291 414
57 414
3 3 23 0 0 0 0 62 61 0 0 4
297 213
291 213
291 359
298 359
4 0 24 0 0 0 0 61 0 0 211 3
322 383
322 430
281 430
4 1 24 0 0 0 0 62 2 0 0 5
321 237
321 273
281 273
281 475
56 475
1 1 100 0 0 4224 0 57 3 0 0 2
82 314
60 314
3 2 101 0 0 4224 0 58 61 0 0 2
276 341
298 341
5 2 102 0 0 12416 0 62 60 0 0 6
351 213
374 213
374 95
136 95
136 168
164 168
2 3 103 0 0 4224 0 56 60 0 0 2
123 177
164 177
3 1 104 0 0 8320 0 59 58 0 0 4
217 305
223 305
223 332
230 332
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
