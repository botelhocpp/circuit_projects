CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 110 30 120 10
125 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
293 176 406 273
9437202 0
0
6 Title:
5 Name:
0
0
0
32
5 4049~
219 707 648 0 2 22
0 3 4
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
8885 0 0
2
45462.5 0
0
7 Ground~
168 756 680 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3780 0 0
2
45462.4 0
0
4 4076
219 805 604 0 22 29
0 12 11 10 9 2 2 2 2 4
2 5 6 7 8 0 0 0 0 0
1 1 1
0
0 0 4848 0
4 4076
-14 -60 14 -52
2 U5
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 14 10 9 2 1 7
15 3 4 5 6 11 12 13 14 10
9 2 1 7 15 3 4 5 6 0
65 0 0 0 0 0 0 0
1 U
9265 0 0
2
45462.4 0
0
14 NO PushButton~
191 517 309 0 2 5
0 18 13
0
0 0 4720 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9442 0 0
2
5.90128e-315 5.32571e-315
0
14 NO PushButton~
191 516 354 0 2 5
0 17 13
0
0 0 4720 0
0
2 S3
-6 -20 8 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9424 0 0
2
5.90128e-315 5.30499e-315
0
14 NO PushButton~
191 517 217 0 2 5
0 20 13
0
0 0 4720 0
0
2 SF
-7 -21 7 -13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9968 0 0
2
5.90128e-315 5.26354e-315
0
14 NO PushButton~
191 517 264 0 2 5
0 19 13
0
0 0 4720 0
0
2 SB
-8 -20 6 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9281 0 0
2
5.90128e-315 0
0
14 NO PushButton~
191 455 308 0 2 5
0 18 14
0
0 0 4720 0
0
2 S6
-8 -20 6 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8464 0 0
2
5.90128e-315 5.32571e-315
0
14 NO PushButton~
191 455 263 0 2 5
0 19 14
0
0 0 4720 0
0
2 SA
-8 -20 6 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7168 0 0
2
5.90128e-315 5.30499e-315
0
14 NO PushButton~
191 455 216 0 2 5
0 20 14
0
0 0 4720 0
0
2 SE
-7 -21 7 -13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3171 0 0
2
5.90128e-315 5.26354e-315
0
14 NO PushButton~
191 454 353 0 2 5
0 17 14
0
0 0 4720 0
0
2 S2
-6 -20 8 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4139 0 0
2
5.90128e-315 0
0
14 NO PushButton~
191 386 353 0 2 5
0 17 15
0
0 0 4720 0
2 S1
-7 -20 7 -12
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 -1 0
1 S
6435 0 0
2
5.90128e-315 5.32571e-315
0
14 NO PushButton~
191 387 308 0 2 5
0 18 15
0
0 0 4720 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5283 0 0
2
5.90128e-315 5.30499e-315
0
14 NO PushButton~
191 387 263 0 2 5
0 19 15
0
0 0 4720 0
0
2 S9
-8 -20 6 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6874 0 0
2
5.90128e-315 5.26354e-315
0
14 NO PushButton~
191 387 216 0 2 5
0 20 15
0
0 0 4720 0
0
2 SD
-7 -21 7 -13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5305 0 0
2
5.90128e-315 0
0
14 NO PushButton~
191 308 354 0 2 5
0 17 16
0
0 0 4720 0
0
2 S0
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
34 0 0
2
5.90128e-315 0
0
14 NO PushButton~
191 309 309 0 2 5
0 18 16
0
0 0 4720 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
969 0 0
2
5.90128e-315 0
0
14 NO PushButton~
191 309 264 0 2 5
0 19 16
0
0 0 4720 0
0
2 S8
-8 -20 6 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8402 0 0
2
5.90128e-315 0
0
14 NO PushButton~
191 309 217 0 2 5
0 20 16
0
0 0 4720 0
0
2 SC
-7 -21 7 -13
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3751 0 0
2
5.90128e-315 0
0
7 Ground~
168 140 679 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4292 0 0
2
45462.4 0
0
7 Ground~
168 679 407 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6118 0 0
2
45462.4 1
0
12 Hex Display~
7 867 528 0 18 19
10 5 6 7 8 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
34 0 0
2
45462.4 2
0
7 74LS293
154 190 578 0 8 17
0 2 2 23 9 12 11 10 9
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U4
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
6357 0 0
2
45462.4 3
0
7 74LS139
118 191 469 0 14 29
0 10 9 2 24 25 26 13 14 15
16 27 28 29 30
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
319 0 0
2
45462.4 4
0
7 74LS153
119 598 426 0 14 29
0 20 19 18 17 12 11 31 32 33
34 2 35 3 36
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
3976 0 0
2
45462.4 5
0
5 4081~
219 112 587 0 3 22
0 22 3 23
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
7634 0 0
2
45462.4 6
0
7 Pulser~
4 37 587 0 10 12
0 37 38 22 39 0 0 10 10 1
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
523 0 0
2
45462.4 7
0
2 +V
167 202 146 0 1 3
0 21
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6748 0 0
2
45462.4 8
0
9 Resistor~
219 147 216 0 4 5
0 17 21 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6901 0 0
2
45462.4 9
0
9 Resistor~
219 185 216 0 4 5
0 18 21 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
842 0 0
2
45462.4 10
0
9 Resistor~
219 219 217 0 4 5
0 19 21 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3277 0 0
2
45462.4 11
0
9 Resistor~
219 254 217 0 4 5
0 20 21 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4212 0 0
2
45462.4 12
0
67
1 0 3 0 0 4096 0 1 0 0 59 2
692 648
657 648
2 9 4 0 0 4224 0 1 3 0 0 4
728 648
754 648
754 649
773 649
0 1 2 0 0 8192 0 0 2 7 0 3
757 658
756 658
756 674
5 0 2 0 0 0 0 3 0 0 5 3
767 613
756 613
756 622
6 0 2 0 0 0 0 3 0 0 7 3
767 622
756 622
756 631
8 0 2 0 0 0 0 3 0 0 7 2
767 640
756 640
7 10 2 0 0 8208 0 3 3 0 0 4
767 631
757 631
757 658
773 658
1 11 5 0 0 4224 0 22 3 0 0 3
876 552
876 595
837 595
12 2 6 0 0 8320 0 3 22 0 0 3
837 586
870 586
870 552
13 3 7 0 0 4224 0 3 22 0 0 3
837 577
864 577
864 552
14 4 8 0 0 4224 0 3 22 0 0 3
837 568
858 568
858 552
8 0 9 0 0 4096 0 23 0 0 22 2
222 596
232 596
0 7 10 0 0 4096 0 0 23 20 0 2
242 587
222 587
0 6 11 0 0 4224 0 0 23 61 0 2
526 578
222 578
1 5 12 0 0 12416 0 3 23 0 0 4
773 568
516 568
516 569
222 569
7 2 13 0 0 4224 0 24 5 0 0 3
229 442
499 442
499 362
8 2 14 0 0 4224 0 24 11 0 0 3
229 451
437 451
437 361
9 2 15 0 0 4224 0 24 12 0 0 3
229 460
369 460
369 361
10 2 16 0 0 8320 0 24 16 0 0 3
229 469
291 469
291 362
3 1 10 0 0 4224 0 3 24 0 0 8
773 586
242 586
242 587
240 587
240 527
119 527
119 451
159 451
0 3 2 0 0 4096 0 0 24 25 0 3
140 569
140 469
153 469
0 2 9 0 0 8192 0 0 24 23 0 5
232 596
232 535
129 535
129 460
159 460
4 4 9 0 0 20608 0 23 3 0 0 6
152 596
131 596
131 650
232 650
232 595
773 595
2 0 2 0 0 0 0 23 0 0 25 2
158 578
140 578
1 1 2 0 0 8320 0 23 20 0 0 3
158 569
140 569
140 673
1 0 17 0 0 12288 0 5 0 0 27 4
533 362
558 362
558 376
485 376
1 0 17 0 0 0 0 11 0 0 28 4
471 361
485 361
485 376
421 376
1 0 17 0 0 12288 0 12 0 0 50 4
403 361
421 361
421 376
343 376
1 0 18 0 0 12288 0 4 0 0 30 4
534 317
558 317
558 327
484 327
1 0 18 0 0 0 0 8 0 0 31 4
472 316
484 316
484 327
421 327
1 0 18 0 0 12288 0 13 0 0 51 4
404 316
421 316
421 327
343 327
1 0 19 0 0 12288 0 7 0 0 33 4
534 272
558 272
558 284
484 284
1 0 19 0 0 0 0 9 0 0 34 4
472 271
484 271
484 284
421 284
1 0 19 0 0 12288 0 14 0 0 52 4
404 271
421 271
421 284
343 284
1 0 20 0 0 12288 0 6 0 0 36 4
534 225
558 225
558 239
484 239
1 0 20 0 0 0 0 10 0 0 37 4
472 224
484 224
484 239
421 239
1 0 20 0 0 12288 0 15 0 0 53 4
404 224
421 224
421 239
343 239
2 2 13 0 0 0 0 4 5 0 0 3
500 317
499 317
499 362
2 2 13 0 0 0 0 7 4 0 0 2
500 272
500 317
2 2 13 0 0 0 0 6 7 0 0 2
500 225
500 272
2 2 14 0 0 0 0 10 9 0 0 2
438 224
438 271
2 2 14 0 0 0 0 8 9 0 0 2
438 316
438 271
2 2 14 0 0 0 0 11 8 0 0 3
437 361
438 361
438 316
2 2 15 0 0 0 0 12 13 0 0 3
369 361
370 361
370 316
2 2 15 0 0 0 0 14 13 0 0 2
370 271
370 316
2 2 15 0 0 0 0 15 14 0 0 2
370 224
370 271
2 2 16 0 0 0 0 17 16 0 0 3
292 317
291 317
291 362
2 2 16 0 0 0 0 18 17 0 0 2
292 272
292 317
2 2 16 0 0 0 0 19 18 0 0 2
292 225
292 272
1 0 17 0 0 12288 0 16 0 0 67 4
325 362
343 362
343 376
147 376
1 0 18 0 0 12288 0 17 0 0 66 4
326 317
343 317
343 327
185 327
1 0 19 0 0 12288 0 18 0 0 58 4
326 272
343 272
343 284
219 284
1 0 20 0 0 12288 0 19 0 0 65 4
326 225
343 225
343 239
254 239
2 0 21 0 0 4096 0 31 0 0 55 2
219 199
219 173
0 2 21 0 0 4096 0 0 32 57 0 3
201 173
254 173
254 199
2 0 21 0 0 0 0 30 0 0 57 2
185 198
185 173
2 1 21 0 0 8320 0 29 28 0 0 4
147 198
147 173
202 173
202 155
2 1 19 0 0 4224 0 25 31 0 0 3
566 399
219 399
219 235
13 2 3 0 0 12416 0 25 26 0 0 6
630 408
657 408
657 658
62 658
62 596
88 596
11 1 2 0 0 0 0 25 21 0 0 3
636 390
679 390
679 401
6 2 11 0 0 0 0 25 3 0 0 6
566 435
526 435
526 578
526 578
526 577
773 577
5 0 12 0 0 0 0 25 0 0 15 3
566 426
516 426
516 569
3 1 22 0 0 4224 0 27 26 0 0 2
61 578
88 578
3 3 23 0 0 4224 0 26 23 0 0 2
133 587
152 587
1 1 20 0 0 8320 0 32 25 0 0 3
254 235
254 390
566 390
3 1 18 0 0 4224 0 25 30 0 0 3
566 408
185 408
185 234
1 4 17 0 0 8320 0 29 25 0 0 3
147 234
147 417
566 417
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
