CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
125 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
293 176 406 273
9437202 0
0
6 Title:
5 Name:
0
0
0
27
14 NO PushButton~
191 426 287 0 2 5
0 7 4
0
0 0 4720 0
0
4 SAST
-13 -20 15 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4129 0 0
2
45462.5 2
0
14 NO PushButton~
191 506 286 0 2 5
0 6 5
0
0 0 4720 0
0
2 S0
-9 -20 5 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6278 0 0
2
45462.5 1
0
14 NO PushButton~
191 575 288 0 2 5
0 7 3
0
0 0 4720 0
0
4 SHAS
-12 -20 16 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3482 0 0
2
45462.5 0
0
14 NO PushButton~
191 505 216 0 2 5
0 7 5
0
0 0 4720 0
0
2 S8
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8323 0 0
2
45462.5 2
0
14 NO PushButton~
191 426 217 0 2 5
0 9 3
0
0 0 4720 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3984 0 0
2
45462.5 1
0
14 NO PushButton~
191 577 216 0 2 5
0 7 8
0
0 0 4720 0
2 S1
-7 -20 7 -12
2 S9
-7 -19 7 -11
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 -1 0
1 S
7622 0 0
2
45462.5 0
0
14 NO PushButton~
191 576 156 0 2 5
0 9 4
0
0 0 4720 0
0
2 S6
-8 -20 6 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
816 0 0
2
45462.5 2
0
14 NO PushButton~
191 504 155 0 2 5
0 9 8
0
0 0 4720 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4656 0 0
2
45462.5 1
0
14 NO PushButton~
191 426 157 0 2 5
0 9 5
0
0 0 4720 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6356 0 0
2
45462.5 0
0
14 NO PushButton~
191 425 90 0 2 5
0 6 8
0
0 0 4720 0
0
2 S1
-8 -20 6 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7479 0 0
2
45462.5 6
0
14 NO PushButton~
191 502 89 0 2 5
0 6 4
0
0 0 4720 0
0
2 S2
-8 -20 6 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5690 0 0
2
45462.5 5
0
14 NO PushButton~
191 573 89 0 2 5
0 6 3
0
0 0 4720 0
0
2 S3
-8 -19 6 -11
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5617 0 0
2
45462.5 4
0
5 4049~
219 707 648 0 2 22
0 11 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
3903 0 0
2
5.90128e-315 0
0
7 Ground~
168 756 680 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4452 0 0
2
5.90128e-315 0
0
4 4076
219 805 604 0 22 29
0 20 19 18 17 2 2 2 2 12
2 13 14 15 16 0 0 0 0 0
1 0 1
0
0 0 4848 0
4 4076
-14 -60 14 -52
2 U5
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 14 10 9 2 1 7
15 3 4 5 6 11 12 13 14 10
9 2 1 7 15 3 4 5 6 0
65 0 0 0 1 0 0 0
1 U
6282 0 0
2
5.90128e-315 0
0
7 Ground~
168 140 679 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7187 0 0
2
5.90128e-315 0
0
7 Ground~
168 679 407 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6866 0 0
2
5.90128e-315 5.26354e-315
0
12 Hex Display~
7 867 528 0 18 19
10 13 14 15 16 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7670 0 0
2
5.90128e-315 5.30499e-315
0
7 74LS293
154 190 578 0 8 17
0 2 2 22 17 20 19 18 17
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U4
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
951 0 0
2
5.90128e-315 5.32571e-315
0
7 74LS139
118 191 469 0 14 29
0 18 17 2 23 24 25 3 4 8
5 26 27 28 29
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
9536 0 0
2
5.90128e-315 5.34643e-315
0
7 74LS153
119 598 426 0 14 29
0 30 7 9 6 20 19 31 32 33
34 2 35 11 36
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
5495 0 0
2
5.90128e-315 5.3568e-315
0
5 4081~
219 112 587 0 3 22
0 21 11 22
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
8152 0 0
2
5.90128e-315 5.36716e-315
0
7 Pulser~
4 37 587 0 10 12
0 37 38 21 39 0 0 10 10 7
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6223 0 0
2
5.90128e-315 5.37752e-315
0
2 +V
167 179 36 0 1 3
0 10
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5441 0 0
2
5.90128e-315 5.38788e-315
0
9 Resistor~
219 140 74 0 4 5
0 7 10 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3189 0 0
2
5.90128e-315 5.39306e-315
0
9 Resistor~
219 179 73 0 4 5
0 9 10 0 1
0
0 0 880 90
3 10k
5 -1 26 7
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8460 0 0
2
5.90128e-315 5.39824e-315
0
9 Resistor~
219 216 75 0 4 5
0 6 10 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5179 0 0
2
5.90128e-315 5.40342e-315
0
57
0 2 3 0 0 4096 0 0 3 19 0 3
283 334
558 334
558 296
0 2 4 0 0 4096 0 0 1 20 0 3
276 327
409 327
409 295
0 2 5 0 0 4096 0 0 2 15 0 3
260 319
489 319
489 294
1 0 6 0 0 12288 0 2 0 0 30 4
523 294
543 294
543 312
216 312
0 1 7 0 0 4096 0 0 3 6 0 4
460 306
609 306
609 296
592 296
1 0 7 0 0 12288 0 1 0 0 28 4
443 295
460 295
460 306
140 306
0 2 8 0 0 4096 0 0 6 21 0 3
268 261
560 261
560 224
0 2 5 0 0 0 0 0 4 15 0 3
260 255
488 255
488 224
0 1 7 0 0 0 0 0 6 10 0 4
543 248
608 248
608 224
594 224
1 0 7 0 0 12288 0 4 0 0 28 4
522 224
543 224
543 248
140 248
0 2 3 0 0 0 0 0 5 19 0 3
283 242
409 242
409 225
1 0 9 0 0 12288 0 5 0 0 29 4
443 225
459 225
459 235
179 235
0 2 4 0 0 4096 0 0 7 20 0 3
276 194
559 194
559 164
0 2 8 0 0 0 0 0 8 21 0 3
268 188
487 188
487 163
10 2 5 0 0 8320 0 20 9 0 0 5
229 469
260 469
260 181
409 181
409 165
0 1 9 0 0 0 0 0 7 17 0 4
543 173
608 173
608 164
593 164
0 1 9 0 0 0 0 0 8 18 0 4
459 173
543 173
543 163
521 163
1 0 9 0 0 0 0 9 0 0 29 4
443 165
459 165
459 174
179 174
7 2 3 0 0 8320 0 20 12 0 0 5
229 442
283 442
283 130
556 130
556 97
8 2 4 0 0 8320 0 20 11 0 0 5
229 451
276 451
276 125
485 125
485 97
9 2 8 0 0 8320 0 20 10 0 0 5
229 460
268 460
268 118
408 118
408 98
0 0 6 0 0 0 0 0 0 24 30 2
459 110
216 110
1 0 6 0 0 0 0 11 0 0 24 3
519 97
543 97
543 110
1 1 6 0 0 0 0 10 12 0 0 6
442 98
459 98
459 110
609 110
609 97
590 97
2 2 10 0 0 8192 0 26 27 0 0 3
179 55
179 57
216 57
2 2 10 0 0 8320 0 26 25 0 0 3
179 55
179 56
140 56
1 2 10 0 0 0 0 24 26 0 0 2
179 45
179 55
2 1 7 0 0 4224 0 21 25 0 0 3
566 399
140 399
140 92
3 1 9 0 0 4224 0 21 26 0 0 3
566 408
179 408
179 91
1 4 6 0 0 8320 0 27 21 0 0 3
216 93
216 417
566 417
1 0 11 0 0 4096 0 13 0 0 52 2
692 648
657 648
2 9 12 0 0 4224 0 13 15 0 0 4
728 648
754 648
754 649
773 649
0 1 2 0 0 8192 0 0 14 37 0 3
757 658
756 658
756 674
5 0 2 0 0 0 0 15 0 0 35 3
767 613
756 613
756 622
6 0 2 0 0 0 0 15 0 0 37 3
767 622
756 622
756 631
8 0 2 0 0 0 0 15 0 0 37 2
767 640
756 640
7 10 2 0 0 8192 0 15 15 0 0 4
767 631
757 631
757 658
773 658
1 11 13 0 0 4224 0 18 15 0 0 3
876 552
876 595
837 595
12 2 14 0 0 8320 0 15 18 0 0 3
837 586
870 586
870 552
13 3 15 0 0 4224 0 15 18 0 0 3
837 577
864 577
864 552
14 4 16 0 0 4224 0 15 18 0 0 3
837 568
858 568
858 552
8 0 17 0 0 4096 0 19 0 0 48 2
222 596
232 596
0 7 18 0 0 4096 0 0 19 46 0 2
242 587
222 587
0 6 19 0 0 4224 0 0 19 54 0 2
526 578
222 578
1 5 20 0 0 12416 0 15 19 0 0 4
773 568
516 568
516 569
222 569
3 1 18 0 0 4224 0 15 20 0 0 8
773 586
242 586
242 587
240 587
240 527
119 527
119 451
159 451
0 3 2 0 0 4096 0 0 20 51 0 3
140 569
140 469
153 469
0 2 17 0 0 8192 0 0 20 49 0 5
232 596
232 535
129 535
129 460
159 460
4 4 17 0 0 20608 0 19 15 0 0 6
152 596
131 596
131 650
232 650
232 595
773 595
2 0 2 0 0 0 0 19 0 0 51 2
158 578
140 578
1 1 2 0 0 8320 0 19 16 0 0 3
158 569
140 569
140 673
13 2 11 0 0 12416 0 21 22 0 0 6
630 408
657 408
657 658
62 658
62 596
88 596
11 1 2 0 0 0 0 21 17 0 0 3
636 390
679 390
679 401
6 2 19 0 0 0 0 21 15 0 0 6
566 435
526 435
526 578
526 578
526 577
773 577
5 0 20 0 0 0 0 21 0 0 45 3
566 426
516 426
516 569
3 1 21 0 0 4224 0 23 22 0 0 2
61 578
88 578
3 3 22 0 0 4224 0 22 19 0 0 2
133 587
152 587
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
