CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 180 30 150 10
133 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
301 176 414 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
7 Ground~
168 212 614 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8809 0 0
2
5.90128e-315 0
0
7 Ground~
168 679 407 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5993 0 0
2
5.90128e-315 0
0
12 Hex Display~
7 766 531 0 18 19
10 7 11 9 10 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8654 0 0
2
5.90128e-315 0
0
7 Ground~
168 337 499 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7223 0 0
2
5.90128e-315 0
0
7 74LS293
154 254 578 0 8 17
0 2 2 13 7 10 9 11 7
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U4
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
3641 0 0
2
5.90128e-315 0
0
7 74LS139
118 386 486 0 14 29
0 11 7 2 19 20 21 6 5 4
3 22 23 24 25
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
3104 0 0
2
5.90128e-315 0
0
7 74LS153
119 598 426 0 14 29
0 6 15 16 17 10 9 26 27 28
29 2 30 8 31
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
3296 0 0
2
5.90128e-315 0
0
5 4081~
219 162 587 0 3 22
0 12 8 13
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
8534 0 0
2
5.90128e-315 0
0
7 Pulser~
4 59 587 0 10 12
0 32 33 12 34 0 0 10 10 3
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
949 0 0
2
5.90128e-315 0
0
2 +V
167 359 196 0 1 3
0 18
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3371 0 0
2
5.90128e-315 0
0
11 4x4 Switch~
193 473 313 0 11 17
0 6 15 16 17 6 3 4 5 0
4 19
0
0 0 4720 0
0
3 SW1
-17 -42 4 -34
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
2 SW
7311 0 0
2
5.90128e-315 0
0
9 Resistor~
219 314 262 0 4 5
0 17 18 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
5.90128e-315 0
0
9 Resistor~
219 343 264 0 4 5
0 16 18 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3526 0 0
2
5.90128e-315 0
0
9 Resistor~
219 374 264 0 4 5
0 15 18 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4129 0 0
2
5.90128e-315 0
0
9 Resistor~
219 403 263 0 4 5
0 6 18 0 1
0
0 0 880 90
3 10k
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6278 0 0
2
5.90128e-315 0
0
32
10 6 3 0 0 8320 0 6 11 0 0 3
424 486
451 486
451 364
9 7 4 0 0 8320 0 6 11 0 0 3
424 477
466 477
466 364
8 8 5 0 0 8320 0 6 11 0 0 3
424 468
480 468
480 364
7 5 6 0 0 8320 0 6 11 0 0 3
424 459
495 459
495 364
0 1 2 0 0 4096 0 0 1 6 0 2
212 576
212 608
1 2 2 0 0 0 0 5 5 0 0 4
222 569
212 569
212 578
222 578
0 4 7 0 0 8192 0 0 5 12 0 5
325 596
325 636
191 636
191 596
216 596
13 2 8 0 0 12416 0 7 8 0 0 6
630 408
657 408
657 658
110 658
110 596
138 596
11 1 2 0 0 4224 0 7 2 0 0 3
636 390
679 390
679 401
6 0 9 0 0 8192 0 7 0 0 14 3
566 435
526 435
526 578
5 0 10 0 0 8192 0 7 0 0 15 3
566 426
517 426
517 569
0 1 7 0 0 4224 0 0 3 18 0 3
325 596
775 596
775 555
2 0 11 0 0 8320 0 3 0 0 17 3
769 555
769 587
316 587
6 3 9 0 0 4224 0 5 3 0 0 3
286 578
763 578
763 555
4 5 10 0 0 8320 0 3 5 0 0 3
757 555
757 569
286 569
3 1 2 0 0 0 0 6 4 0 0 3
348 486
337 486
337 493
7 1 11 0 0 0 0 5 6 0 0 4
286 587
319 587
319 468
354 468
2 8 7 0 0 0 0 6 5 0 0 4
354 477
325 477
325 596
286 596
3 1 12 0 0 4224 0 9 8 0 0 2
83 578
138 578
3 3 13 0 0 4224 0 8 5 0 0 2
183 587
216 587
0 1 6 0 0 8320 14 0 7 32 0 3
403 291
403 390
566 390
0 2 15 0 0 8320 0 0 7 31 0 3
375 306
375 399
566 399
3 0 16 0 0 4224 0 7 0 0 30 3
566 408
343 408
343 319
0 4 17 0 0 8320 0 0 7 29 0 3
314 335
314 417
566 417
1 0 18 0 0 4224 0 10 0 0 27 2
359 205
359 238
0 2 18 0 0 0 0 0 15 27 0 3
374 238
403 238
403 245
0 2 18 0 0 0 0 0 14 28 0 3
343 238
374 238
374 246
2 2 18 0 0 0 0 12 13 0 0 4
314 244
314 238
343 238
343 246
4 1 17 0 0 0 0 11 12 0 0 3
422 335
314 335
314 280
1 3 16 0 0 0 0 13 11 0 0 3
343 282
343 320
422 320
2 1 15 0 0 0 0 11 14 0 0 3
422 306
374 306
374 282
1 1 6 0 0 0 14 11 15 0 0 3
422 291
403 291
403 281
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
